* C:\FOSSEE\eSim\library\SubcircuitLibrary\astable_multivibrator\astable_multivibrator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/05/22 22:03:57

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_C1-Pad1_ Net-_R1-Pad2_ 10k		
R3  Net-_R3-Pad1_ Net-_R1-Pad2_ 1k		
R4  GND Net-_R3-Pad1_ 10k		
C1  Net-_C1-Pad1_ GND 0.01u		
v1  Net-_X1-Pad7_ GND 5V		
X1  Net-_R2-Pad1_ Net-_C1-Pad1_ Net-_R3-Pad1_ GND Net-_R2-Pad2_ Net-_R1-Pad2_ Net-_X1-Pad7_ ? lm_741		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 1k		
U1  Net-_R1-Pad2_ PORT		

.end
